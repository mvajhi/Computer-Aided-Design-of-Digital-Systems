module Counter4bit (
    input clk,
    input rst,
);
        
endmodule