module Read_Controller_Filter(
    input co_Filter,
    input av_input,
    input Filter_size,
    input write_pointer,
    input read_pointer,
    
    output write_en_src_pad,
    output write_counter_en,
    output end_of_filter,
    output av_filter
);

endmodule