module dp #(
    parameter IFMAP_BUFFER_WIDTH = 18,
) (
    input clk,
    input rst,
    input start,
);

endmodule