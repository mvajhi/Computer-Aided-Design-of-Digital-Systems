module ReadAddressGeneratorFilter (
    input clk,
    input rst,
);

endmodule